bplist00�SURL_efile:///Users/manuel/Library/Messages/Attachments/eb/11/B3BB95E8-E13A-4155-B97D-25E9E0C4A6DD/alarm.sv                            w